
module short (a, a);
    inout a;
endmodule
