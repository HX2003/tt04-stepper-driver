
module short (.ioa(a), .iob(a));
    inout a;
endmodule
